<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,120.8,-89.2</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>12,-12.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>12,-15.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>23,-12</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_SMALL_INVERTER</type>
<position>23,-14.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>36,-12.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>36,-18</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>36,-24</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>36,-29.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>50,-17</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>53.5,-17</position>
<input>
<ID>N_in2</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>57,-17</position>
<input>
<ID>N_in2</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>60.5,-17</position>
<input>
<ID>N_in2</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-12.5,21,-12.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>19 2</intersection>
<intersection>21 6</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>19,-30.5,19,-12.5</points>
<intersection>-30.5 3</intersection>
<intersection>-17 5</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>19,-30.5,33,-30.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>19 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>19,-17,33,-17</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>19 2</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>21,-12.5,21,-12</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-15.5,21,-15.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>21 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21,-28.5,21,-14.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-28.5 6</intersection>
<intersection>-23 4</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>21,-23,33,-23</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>21 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>21,-28.5,33,-28.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>21 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-12,29,-11.5</points>
<intersection>-12 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-11.5,33,-11.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection>
<intersection>31 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-12,29,-12</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>31,-25,31,-11.5</points>
<intersection>-25 5</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>31,-25,33,-25</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>31 4</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-19,29,-13.5</points>
<intersection>-19 4</intersection>
<intersection>-14.5 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-13.5,33,-13.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-14.5,29,-14.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>29,-19,33,-19</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-17,44,-12.5</points>
<intersection>-17 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-17,49,-17</points>
<connection>
<GID>18</GID>
<name>N_in0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-12.5,44,-12.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-19,53.5,-19</points>
<intersection>39 2</intersection>
<intersection>53.5 3</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>39,-19,39,-18</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>-19 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>53.5,-19,53.5,-18</points>
<connection>
<GID>20</GID>
<name>N_in2</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-24,57,-18</points>
<connection>
<GID>22</GID>
<name>N_in2</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-24,57,-24</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-29.5,60.5,-18</points>
<connection>
<GID>24</GID>
<name>N_in2</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-29.5,60.5,-29.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,120.8,-89.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,120.8,-89.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,120.8,-89.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,120.8,-89.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,120.8,-89.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,120.8,-89.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,120.8,-89.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,120.8,-89.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,120.8,-89.2</PageViewport></page 9></circuit>