<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>29,-17.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>29,-26</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>44,-17</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND2</type>
<position>43.5,-26</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>35.5,-17.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>34.5,-26</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_SMALL_INVERTER</type>
<position>51,-16.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_SMALL_INVERTER</type>
<position>50.5,-26</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>17,-29.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>17,-27</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>57.5,-22</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AE_SMALL_INVERTER</type>
<position>21.5,-20.5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-17.5,33.5,-17.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-17.5,39,-16</points>
<intersection>-17.5 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-16,41,-16</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-17.5,39,-17.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32,-26,32.5,-26</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-27,38.5,-26</points>
<intersection>-27 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-27,40.5,-27</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-26,38.5,-26</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,-16.5,49,-16.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>47 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>47,-17,47,-16.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-22,49,-20</points>
<intersection>-22 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-22,49,-22</points>
<intersection>40.5 3</intersection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-20,54.5,-20</points>
<intersection>49 0</intersection>
<intersection>54.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40.5,-25,40.5,-22</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-22 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>54.5,-20,54.5,-16.5</points>
<intersection>-20 2</intersection>
<intersection>-16.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>53,-16.5,54.5,-16.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>54.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-26,48.5,-26</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-21,53.5,-21</points>
<intersection>41 3</intersection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41,-21,41,-18</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-21 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-26,53.5,-21</points>
<intersection>-26 15</intersection>
<intersection>-22 10</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>53.5,-22,56.5,-22</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>53.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>52.5,-26,53.5,-26</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>53.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-29.5,24,-18.5</points>
<intersection>-29.5 3</intersection>
<intersection>-25 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-18.5,26,-18.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-25,26,-25</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>19,-29.5,24,-29.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-18.5,21.5,-14.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-14.5,26,-14.5</points>
<intersection>21.5 0</intersection>
<intersection>26 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>26,-16.5,26,-14.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-27,26,-27</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>21.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21.5,-27,21.5,-22.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport></page 1>
<page 2>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport></page 2>
<page 3>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport></page 3>
<page 4>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport></page 4>
<page 5>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport></page 5>
<page 6>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport></page 6>
<page 7>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport></page 7>
<page 8>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport></page 8>
<page 9>
<PageViewport>0,2.6526e-006,120.8,-89.2</PageViewport></page 9></circuit>